module message #(
	parameter LEN = 8,		
)(
	input raw_i,
);

endmodule

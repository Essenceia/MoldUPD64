module message_block #(
	parameter LEN = 8,		
)(
	input raw_i,
);

endmodule
